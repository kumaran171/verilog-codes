module xnor_gate_struct(output Y,input A,B);
   xnor g1(Y,A,B);
endmodule