module nor_gate_struct(output Y, input A,B);
    nor g1(Y,A,B);
endmodule