module xor_gate_struc(output Y, input A, input B);
  xor g1(Y, A, B);
endmodule