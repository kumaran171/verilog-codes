module or_gate_structural(output Y, input A, input B);
    or g1(Y, A, B);
endmodule