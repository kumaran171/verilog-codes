$date
	Tue May 27 15:44:21 2025
$end
$version
	Icarus Verilog
$end
$timescale
	1s
$end
$scope module tb_not_dat $end
$var wire 1 ! y $end
$var reg 1 " a $end
$scope module uut $end
$var wire 1 # A $end
$var wire 1 ! Y $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0#
0"
1!
$end
#10
0!
1"
1#
#20
