module or_gate_dataflow(output Y, input A, input B);
     assign Y=A | B;
endmodule