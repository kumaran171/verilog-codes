module not_gate_struct(output Y,input A);
   not g1(Y,A);
endmodule