module nand_gate_struc(output Y,input A,B);
  nand g1(Y,A,B);
endmodule