module xor_data(output Y, input A,B);
  assign Y=A ^ B;
endmodule