module tb_8_3_enc_s;
  reg [7:0] d;
  wire [2:0] a;
  enco_8_3_s uut(.d(d),.a(a));
  initial begin
    $dumpfile("z16.vcd");
    $dumpvars(0,tb_8_3_enc_s);
    $display("D7 D6 D5 D4 D3 D2 D1 D0 | A2 A1 A0");
    $monitor("%b %b %b %b %b %b %b %b| %b %b %b",d[7],d[6],d[5],d[4],d[3],d[2],d[1],d[0],a[2],a[1],a[0]);
    d[7]=1;d[6]=0;d[5]=0;d[4]=0;d[3]=0;d[2]=0;d[1]=0;d[0]=0;#10;
    d[7]=0;d[6]=1;d[5]=0;d[4]=0;d[3]=0;d[2]=0;d[1]=0;d[0]=0;#10;
    d[7]=0;d[6]=0;d[5]=1;d[4]=0;d[3]=0;d[2]=0;d[1]=0;d[0]=0;#10;
    d[7]=0;d[6]=0;d[5]=0;d[4]=1;d[3]=0;d[2]=0;d[1]=0;d[0]=0;#10;
    d[7]=0;d[6]=0;d[5]=0;d[4]=0;d[3]=1;d[2]=0;d[1]=0;d[0]=0;#10;
    d[7]=0;d[6]=0;d[5]=0;d[4]=0;d[3]=0;d[2]=1;d[1]=0;d[0]=0;#10;
    d[7]=0;d[6]=0;d[5]=0;d[4]=0;d[3]=0;d[2]=0;d[1]=1;d[0]=0;#10;
    d[7]=0;d[6]=0;d[5]=0;d[4]=0;d[3]=0;d[2]=0;d[1]=0;d[0]=1;#10;
    d[7]=0;d[6]=0;d[5]=0;d[4]=0;d[3]=0;d[2]=0;d[1]=0;d[0]=0;#10;
    $finish;
 end
endmodule






    
    