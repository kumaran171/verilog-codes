module and_gate_data(output Y, input A, input B);
  assign Y=A & B;
endmodule