module not_gate_dat(output Y,input A);
   assign Y=~A;
endmodule