module and_gate_structural(output Y, input A, B);
  and g1(Y, A, B);  
endmodule
